RECT 0.0 -24.87 2.5 24.87 ;
RECT 2.5 -24.49 5.0 24.49 ;
RECT 5.0 -23.85 7.5 23.85 ;
RECT 7.5 -22.91 10.0 22.91 ;
RECT 10.0 -21.65 12.5 21.65 ;
RECT 12.5 -20.0 15.0 20.0 ;
RECT 15.0 -17.85 17.5 17.85 ;
RECT 17.5 -15.0 20.0 15.0 ;
RECT 20.0 -10.9 22.5 10.9 ;
RECT 22.5 -0.0 25.0 0.0 ;
RECT -2.5 -24.87 -0.0 24.87 ;
RECT -5.0 -24.49 -2.5 24.49 ;
RECT -7.5 -23.85 -5.0 23.85 ;
RECT -10.0 -22.91 -7.5 22.91 ;
RECT -12.5 -21.65 -10.0 21.65 ;
RECT -15.0 -20.0 -12.5 20.0 ;
RECT -17.5 -17.85 -15.0 17.85 ;
RECT -20.0 -15.0 -17.5 15.0 ;
RECT -22.5 -10.9 -20.0 10.9 ;
RECT -25.0 -0.0 -22.5 0.0 ;
